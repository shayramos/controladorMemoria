module FIFOFull();


endmodule
