module FIFOEmpty();


endmodule
